module jt900h;

endmodule